package cnt_pkg;
	int test_finished = 0;
	int error_count = 0;
	int correct_count = 0;
	event etrigger;
endpackage : cnt_pkg